module carry_skip_adder
#(
    parameter DATA_WIDTH = 16
)(
    input wire [DATA_WIDTH-1:0] iv_a,
    input wire [DATA_WIDTH-1:0] iv_b,
    input wire i_cin,
    output wire [DATA_WIDTH-1:0] ov_sum,
    output wire o_cout
);

    // WIP



endmodule
