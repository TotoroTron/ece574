module skip_logic
#(
    parameter BLOCK_WIDTH = 4
)(
    input wire [BLOCK_WIDTH-1:0] iv_a,
    input wire [BLOCK_WIDTH-1:0] iv_b,
    input wire i_cin,
    input wire i_rca_cout,
    output wire o_cout
);

    wire [BLOCK_WIDTH-1:0] p;
    wire block_prop;
    
    // WIP!


endmodule
    

